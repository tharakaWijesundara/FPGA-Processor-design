module processorModule (
    
);

alu ALU()
registor_with_inc PC();
    
endmodule