
module ram #(
    parameter DATA_LEN = 16,
    parameter ADDRESS_LEN = 8,
    parameter NO_OF_CORES = 3
)
(
    input clk,
    input read, 
    input write,
    input [ADDRESS_LEN * NO_OF_CORES - 1:0] address,
    input [DATA_LEN * NO_OF_CORES - 1:0] data_in,
    output reg [DATA_LEN * NO_OF_CORES - 1:0] data_out
);
reg [DATA_LEN - 1:0] memory [2 ** ADDRESS_LEN - 1:0];
 initial begin
        memory[0] = 6'd4;
        memory[1] = 12'h3E;
        memory[2] = 6'd36;
        memory[3] = 6'd4;
        memory[4] = 12'h3F;
        memory[5] = 6'd37;
        memory[6] = 6'd14;

		memory[7] = 12'h208;

		memory[8] = 6'd16;
		memory[9] = 12'h388;

		memory[10] = 6'd12;
		memory[11] = 12'h40;

            memory[12] = 12'd58;
            memory[13] = 6'd4;
            memory[14] = 12'd11;
            memory[15] = 12'd39;
            memory[16] = 6'd8;
            memory[17] = 12'd11;
            memory[18] = 6'd4;
            memory[19] = 12'd9;
            memory[20] = 12'd40;
            memory[21] = 6'd8;
            memory[22] = 12'd9;
            memory[23] = 6'd18;
            memory[24] = 6'd38;
            memory[25] = 6'd21;
            memory[26] = 6'd51;
            memory[27] = 6'd38;
            memory[28] = 6'd24;
            memory[29] = 6'd41;
            memory[30] = 6'd33;
            memory[31] = 6'd43;
            memory[32] = 6'd44;
            memory[33] = 6'd4;
            memory[34] = 12'h3D;
            memory[35] = 6'd48;
            memory[36] = 6'd8;
            memory[37] = 12'h3D;
            memory[38] = 6'd46;
            memory[39] = 6'd52;
            memory[40] = 12'h17;
            memory[41] = 6'd42;
            memory[42] = 6'd55;
            memory[43] = 6'd8;
            memory[44] = 12'h3D;
            memory[45] = 6'd4;
            memory[46] = 12'h3C;
            memory[47] = 6'd48;
            memory[48] = 6'd8;
            memory[49] = 12'h3C;
            memory[50] = 6'd45;
            memory[51] = 6'd59;
            memory[52] = 6'd52;
            memory[53] = 12'h17;
            memory[54] = 6'd56;
            memory[55] = 6'd55;
            memory[56] = 6'd8;
            memory[57] = 12'h3C;
            memory[58] = 6'd57;
    end 
 
        initial begin
        memory[60] = 16'd0;
        memory[61] = 16'd0;

		memory[62] = 16'd24;
		memory[63] = 16'd16;
		memory[64] =16'd10;
		memory[65] =16'd38;
		memory[66] =16'd30;
		memory[67] =16'd4;
		memory[68] =16'd19;
		memory[69] =16'd33;
		memory[70] =16'd26;
		memory[71] =16'd5;
		memory[72] =16'd8;
		memory[73] =16'd33;
		memory[74] =16'd41;
		memory[75] =16'd3;
		memory[76] =16'd42;
		memory[77] =16'd40;
		memory[78] =16'd12;
		memory[79] =16'd25;
		memory[80] =16'd40;
		memory[81] =16'd47;
		memory[82] =16'd47;
		memory[83] =16'd46;
		memory[84] =16'd25;
		memory[85] =16'd25;
		memory[86] =16'd24;
		memory[87] =16'd14;
		memory[88] =16'd23;
		memory[89] =16'd16;
		memory[90] =16'd21;
		memory[91] =16'd1;
		memory[92] =16'd23;
		memory[93] =16'd10;
		memory[94] =16'd45;
		memory[95] =16'd42;
		memory[96] =16'd48;
		memory[97] =16'd10;
		memory[98] =16'd26;
		memory[99] =16'd22;
		memory[100] =16'd1;
		memory[101] =16'd32;
		memory[102] =16'd9;
		memory[103] =16'd1;
		memory[104] =16'd4;
		memory[105] =16'd39;
		memory[106] =16'd17;
		memory[107] =16'd26;
		memory[108] =16'd8;
		memory[109] =16'd40;
		memory[110] =16'd38;
		memory[111] =16'd44;
		memory[112] =16'd28;
		memory[113] =16'd7;
		memory[114] =16'd18;
		memory[115] =16'd13;
		memory[116] =16'd47;
		memory[117] =16'd7;
		memory[118] =16'd37;
		memory[119] =16'd13;
		memory[120] =16'd18;
		memory[121] =16'd42;
		memory[122] =16'd11;
		memory[123] =16'd17;
		memory[124] =16'd42;
		memory[125] =16'd6;
		memory[126] =16'd0;
		memory[127] =16'd38;
		memory[128] =16'd24;
		memory[129] =16'd20;
		memory[130] =16'd23;
		memory[131] =16'd34;
		memory[132] =16'd31;
		memory[133] =16'd12;
		memory[134] =16'd12;
		memory[135] =16'd34;
		memory[136] =16'd25;
		memory[137] =16'd6;
		memory[138] =16'd25;
		memory[139] =16'd22;
		memory[140] =16'd2;
		memory[141] =16'd26;
		memory[142] =16'd17;
		memory[143] =16'd0;
		memory[144] =16'd10;
		memory[145] =16'd23;
		memory[146] =16'd31;
		memory[147] =16'd24;
		memory[148] =16'd37;
		memory[149] =16'd5;
		memory[150] =16'd0;
		memory[151] =16'd24;
		memory[152] =16'd47;
		memory[153] =16'd25;
		memory[154] =16'd38;
		memory[155] =16'd44;
		memory[156] =16'd30;
		memory[157] =16'd42;
		memory[158] =16'd35;
		memory[159] =16'd8;
		memory[160] =16'd29;
		memory[161] =16'd3;
		memory[162] =16'd33;
		memory[163] =16'd13;
		memory[164] =16'd30;
		memory[165] =16'd20;
		memory[166] =16'd3;
		memory[167] =16'd48;
		memory[168] =16'd47;
		memory[169] =16'd8;
		memory[170] =16'd19;
		memory[171] =16'd37;
		memory[172] =16'd39;
		memory[173] =16'd35;
		memory[174] =16'd3;
		memory[175] =16'd9;
		memory[176] =16'd45;
		memory[177] =16'd30;
		memory[178] =16'd21;
		memory[179] =16'd6;
		memory[180] =16'd35;
		memory[181] =16'd49;
		memory[182] =16'd26;
		memory[183] =16'd1;
		memory[184] =16'd42;
		memory[185] =16'd43;
		memory[186] =16'd48;
		memory[187] =16'd36;
		memory[188] =16'd9;
		memory[189] =16'd37;
		memory[190] =16'd49;
		memory[191] =16'd16;
		memory[192] =16'd46;
		memory[193] =16'd34;
		memory[194] =16'd20;
		memory[195] =16'd10;
		memory[196] =16'd48;
		memory[197] =16'd47;
		memory[198] =16'd34;
		memory[199] =16'd40;
		memory[200] =16'd41;
		memory[201] =16'd46;
		memory[202] =16'd30;
		memory[203] =16'd23;
		memory[204] =16'd47;
		memory[205] =16'd15;
		memory[206] =16'd24;
		memory[207] =16'd44;
		memory[208] =16'd24;
		memory[209] =16'd40;
		memory[210] =16'd33;
		memory[211] =16'd29;
		memory[212] =16'd40;
		memory[213] =16'd34;
		memory[214] =16'd39;
		memory[215] =16'd44;
		memory[216] =16'd32;
		memory[217] =16'd34;
		memory[218] =16'd47;
		memory[219] =16'd12;
		memory[220] =16'd16;
		memory[221] =16'd8;
		memory[222] =16'd35;
		memory[223] =16'd5;
		memory[224] =16'd15;
		memory[225] =16'd48;
		memory[226] =16'd30;
		memory[227] =16'd38;
		memory[228] =16'd12;
		memory[229] =16'd5;
		memory[230] =16'd31;
		memory[231] =16'd31;
		memory[232] =16'd2;
		memory[233] =16'd46;
		memory[234] =16'd28;
		memory[235] =16'd28;
		memory[236] =16'd25;
		memory[237] =16'd16;
		memory[238] =16'd39;
		memory[239] =16'd24;
		memory[240] =16'd36;
		memory[241] =16'd14;
		memory[242] =16'd24;
		memory[243] =16'd41;
		memory[244] =16'd43;
		memory[245] =16'd28;
		memory[246] =16'd12;
		memory[247] =16'd5;
		memory[248] =16'd18;
		memory[249] =16'd17;
		memory[250] =16'd26;
		memory[251] =16'd21;
		memory[252] =16'd2;
		memory[253] =16'd27;
		memory[254] =16'd36;
		memory[255] =16'd32;
		memory[256] =16'd7;
		memory[257] =16'd49;
		memory[258] =16'd14;
		memory[259] =16'd46;
		memory[260] =16'd49;
		memory[261] =16'd0;
		memory[262] =16'd49;
		memory[263] =16'd40;
		memory[264] =16'd29;
		memory[265] =16'd49;
		memory[266] =16'd12;
		memory[267] =16'd26;
		memory[268] =16'd19;
		memory[269] =16'd3;
		memory[270] =16'd38;
		memory[271] =16'd21;
		memory[272] =16'd10;
		memory[273] =16'd23;
		memory[274] =16'd12;
		memory[275] =16'd38;
		memory[276] =16'd32;
		memory[277] =16'd22;
		memory[278] =16'd43;
		memory[279] =16'd31;
		memory[280] =16'd1;
		memory[281] =16'd20;
		memory[282] =16'd17;
		memory[283] =16'd37;
		memory[284] =16'd6;
		memory[285] =16'd27;
		memory[286] =16'd38;
		memory[287] =16'd48;
		memory[288] =16'd29;
		memory[289] =16'd21;
		memory[290] =16'd9;
		memory[291] =16'd20;
		memory[292] =16'd8;
		memory[293] =16'd14;
		memory[294] =16'd46;
		memory[295] =16'd27;
		memory[296] =16'd3;
		memory[297] =16'd25;
		memory[298] =16'd9;
		memory[299] =16'd33;
		memory[300] =16'd30;
		memory[301] =16'd21;
		memory[302] =16'd34;
		memory[303] =16'd48;
		memory[304] =16'd30;
		memory[305] =16'd13;
		memory[306] =16'd31;
		memory[307] =16'd12;
		memory[308] =16'd21;
		memory[309] =16'd40;
		memory[310] =16'd44;
		memory[311] =16'd20;
		memory[312] =16'd31;
		memory[313] =16'd4;
		memory[314] =16'd16;
		memory[315] =16'd25;
		memory[316] =16'd33;
		memory[317] =16'd18;
		memory[318] =16'd35;
		memory[319] =16'd11;
		memory[320] =16'd8;
		memory[321] =16'd33;
		memory[322] =16'd4;
		memory[323] =16'd19;
		memory[324] =16'd48;
		memory[325] =16'd25;
		memory[326] =16'd7;
		memory[327] =16'd2;
		memory[328] =16'd21;
		memory[329] =16'd37;
		memory[330] =16'd4;
		memory[331] =16'd10;
		memory[332] =16'd18;
		memory[333] =16'd22;
		memory[334] =16'd6;
		memory[335] =16'd33;
		memory[336] =16'd47;
		memory[337] =16'd37;
		memory[338] =16'd46;
		memory[339] =16'd29;
		memory[340] =16'd12;
		memory[341] =16'd15;
		memory[342] =16'd13;
		memory[343] =16'd19;
		memory[344] =16'd6;
		memory[345] =16'd10;
		memory[346] =16'd33;
		memory[347] =16'd14;
		memory[348] =16'd16;
		memory[349] =16'd15;
		memory[350] =16'd44;
		memory[351] =16'd9;
		memory[352] =16'd48;
		memory[353] =16'd31;
		memory[354] =16'd20;
		memory[355] =16'd49;
		memory[356] =16'd43;
		memory[357] =16'd22;
		memory[358] =16'd36;
		memory[359] =16'd28;
		memory[360] =16'd5;
		memory[361] =16'd2;
		memory[362] =16'd44;
		memory[363] =16'd48;
		memory[364] =16'd8;
		memory[365] =16'd17;
		memory[366] =16'd43;
		memory[367] =16'd2;
		memory[368] =16'd9;
		memory[369] =16'd16;
		memory[370] =16'd27;
		memory[371] =16'd6;
		memory[372] =16'd48;
		memory[373] =16'd41;
		memory[374] =16'd10;
		memory[375] =16'd8;
		memory[376] =16'd31;
		memory[377] =16'd38;
		memory[378] =16'd13;
		memory[379] =16'd21;
		memory[380] =16'd12;
		memory[381] =16'd33;
		memory[382] =16'd36;
		memory[383] =16'd4;
		memory[384] =16'd19;
		memory[385] =16'd23;
		memory[386] =16'd20;
		memory[387] =16'd20;
		memory[388] =16'd5;
		memory[389] =16'd8;
		memory[390] =16'd29;
		memory[391] =16'd15;
		memory[392] =16'd43;
		memory[393] =16'd40;
		memory[394] =16'd10;
		memory[395] =16'd8;
		memory[396] =16'd10;
		memory[397] =16'd4;
		memory[398] =16'd10;
		memory[399] =16'd34;
		memory[400] =16'd32;
		memory[401] =16'd29;
		memory[402] =16'd1;
		memory[403] =16'd19;
		memory[404] =16'd41;
		memory[405] =16'd11;
		memory[406] =16'd37;
		memory[407] =16'd18;
		memory[408] =16'd33;
		memory[409] =16'd0;
		memory[410] =16'd43;
		memory[411] =16'd47;
		memory[412] =16'd10;
		memory[413] =16'd46;
		memory[414] =16'd2;
		memory[415] =16'd39;
		memory[416] =16'd27;
		memory[417] =16'd3;
		memory[418] =16'd13;
		memory[419] =16'd32;
		memory[420] =16'd11;
		memory[421] =16'd35;
		memory[422] =16'd22;
		memory[423] =16'd34;
		memory[424] =16'd9;
		memory[425] =16'd27;
		memory[426] =16'd49;
		memory[427] =16'd17;
		memory[428] =16'd35;
		memory[429] =16'd5;
		memory[430] =16'd8;
		memory[431] =16'd28;
		memory[432] =16'd1;
		memory[433] =16'd24;
		memory[434] =16'd24;
		memory[435] =16'd39;
		memory[436] =16'd1;
		memory[437] =16'd37;
		memory[438] =16'd28;
		memory[439] =16'd44;
		memory[440] =16'd29;
		memory[441] =16'd39;
		memory[442] =16'd4;
		memory[443] =16'd16;
		memory[444] =16'd5;
		memory[445] =16'd30;
		memory[446] =16'd18;
		memory[447] =16'd10;
		memory[448] =16'd36;
		memory[449] =16'd7;
		memory[450] =16'd19;
		memory[451] =16'd32;
		memory[452] =16'd44;
		memory[453] =16'd38;
		memory[454] =16'd35;
		memory[455] =16'd16;
		memory[456] =16'd34;
		memory[457] =16'd9;
		memory[458] =16'd42;
		memory[459] =16'd2;
		memory[460] =16'd1;
		memory[461] =16'd28;
		memory[462] =16'd42;
		memory[463] =16'd7;
		memory[464] =16'd40;
		memory[465] =16'd9;
		memory[466] =16'd17;
		memory[467] =16'd22;
		memory[468] =16'd10;
		memory[469] =16'd23;
		memory[470] =16'd4;
		memory[471] =16'd46;
		memory[472] =16'd35;
		memory[473] =16'd11;
		memory[474] =16'd45;
		memory[475] =16'd47;
		memory[476] =16'd6;
		memory[477] =16'd46;
		memory[478] =16'd17;
		memory[479] =16'd45;
		memory[480] =16'd7;
		memory[481] =16'd49;
		memory[482] =16'd37;
		memory[483] =16'd21;
		memory[484] =16'd33;
		memory[485] =16'd44;
		memory[486] =16'd4;
		memory[487] =16'd26;
		memory[488] =16'd24;
		memory[489] =16'd5;
		memory[490] =16'd38;
		memory[491] =16'd42;
		memory[492] =16'd41;
		memory[493] =16'd31;
		memory[494] =16'd1;
		memory[495] =16'd12;
		memory[496] =16'd40;
		memory[497] =16'd20;
		memory[498] =16'd42;
		memory[499] =16'd2;
		memory[500] =16'd15;
		memory[501] =16'd48;
		memory[502] =16'd45;
		memory[503] =16'd18;
		memory[504] =16'd6;
		memory[505] =16'd36;
		memory[506] =16'd35;
		memory[507] =16'd10;
		memory[508] =16'd47;
		memory[509] =16'd21;
		memory[510] =16'd36;
		memory[511] =16'd8;
		memory[512] =16'd32;
		memory[513] =16'd40;
		memory[514] =16'd43;
		memory[515] =16'd0;
		memory[516] =16'd32;
		memory[517] =16'd22;
		memory[518] =16'd47;
		memory[519] =16'd37;

		memory[520] =16'd37;
		memory[521] =16'd13;
		memory[522] =16'd17;
		memory[523] =16'd42;
		memory[524] =16'd26;
		memory[525] =16'd42;
		memory[526] =16'd32;
		memory[527] =16'd3;
		memory[528] =16'd39;
		memory[529] =16'd36;
		memory[530] =16'd35;
		memory[531] =16'd14;
		memory[532] =16'd14;
		memory[533] =16'd45;
		memory[534] =16'd35;
		memory[535] =16'd45;
		memory[536] =16'd27;
		memory[537] =16'd16;
		memory[538] =16'd0;
		memory[539] =16'd27;
		memory[540] =16'd47;
		memory[541] =16'd32;
		memory[542] =16'd30;
		memory[543] =16'd19;
		memory[544] =16'd32;
		memory[545] =16'd48;
		memory[546] =16'd31;
		memory[547] =16'd41;
		memory[548] =16'd48;
		memory[549] =16'd35;
		memory[550] =16'd42;
		memory[551] =16'd28;
		memory[552] =16'd0;
		memory[553] =16'd20;
		memory[554] =16'd15;
		memory[555] =16'd30;
		memory[556] =16'd44;
		memory[557] =16'd0;
		memory[558] =16'd18;
		memory[559] =16'd43;
		memory[560] =16'd1;
		memory[561] =16'd10;
		memory[562] =16'd27;
		memory[563] =16'd33;
		memory[564] =16'd38;
		memory[565] =16'd27;
		memory[566] =16'd26;
		memory[567] =16'd48;
		memory[568] =16'd41;
		memory[569] =16'd10;
		memory[570] =16'd4;
		memory[571] =16'd20;
		memory[572] =16'd7;
		memory[573] =16'd9;
		memory[574] =16'd33;
		memory[575] =16'd10;
		memory[576] =16'd29;
		memory[577] =16'd37;
		memory[578] =16'd20;
		memory[579] =16'd3;
		memory[580] =16'd17;
		memory[581] =16'd15;
		memory[582] =16'd47;
		memory[583] =16'd13;
		memory[584] =16'd27;
		memory[585] =16'd4;
		memory[586] =16'd10;
		memory[587] =16'd5;
		memory[588] =16'd44;
		memory[589] =16'd42;
		memory[590] =16'd3;
		memory[591] =16'd1;
		memory[592] =16'd46;
		memory[593] =16'd30;
		memory[594] =16'd17;
		memory[595] =16'd18;
		memory[596] =16'd10;
		memory[597] =16'd0;
		memory[598] =16'd12;
		memory[599] =16'd6;
		memory[600] =16'd11;
		memory[601] =16'd41;
		memory[602] =16'd41;
		memory[603] =16'd11;
		memory[604] =16'd15;
		memory[605] =16'd35;
		memory[606] =16'd20;
		memory[607] =16'd29;
		memory[608] =16'd3;
		memory[609] =16'd7;
		memory[610] =16'd43;
		memory[611] =16'd34;
		memory[612] =16'd39;
		memory[613] =16'd14;
		memory[614] =16'd24;
		memory[615] =16'd36;
		memory[616] =16'd22;
		memory[617] =16'd9;
		memory[618] =16'd6;
		memory[619] =16'd44;
		memory[620] =16'd46;
		memory[621] =16'd25;
		memory[622] =16'd38;
		memory[623] =16'd46;
		memory[624] =16'd42;
		memory[625] =16'd49;
		memory[626] =16'd4;
		memory[627] =16'd36;
		memory[628] =16'd27;
		memory[629] =16'd42;
		memory[630] =16'd35;
		memory[631] =16'd5;
		memory[632] =16'd41;
		memory[633] =16'd23;
		memory[634] =16'd34;
		memory[635] =16'd47;
		memory[636] =16'd6;
		memory[637] =16'd40;
		memory[638] =16'd1;
		memory[639] =16'd5;
		memory[640] =16'd16;
		memory[641] =16'd27;
		memory[642] =16'd4;
		memory[643] =16'd42;
		memory[644] =16'd25;
		memory[645] =16'd15;
		memory[646] =16'd35;
		memory[647] =16'd29;
		memory[648] =16'd29;
		memory[649] =16'd24;
		memory[650] =16'd40;
		memory[651] =16'd43;
		memory[652] =16'd37;
		memory[653] =16'd43;
		memory[654] =16'd14;
		memory[655] =16'd10;
		memory[656] =16'd30;
		memory[657] =16'd49;
		memory[658] =16'd33;
		memory[659] =16'd20;
		memory[660] =16'd8;
		memory[661] =16'd17;
		memory[662] =16'd34;
		memory[663] =16'd31;
		memory[664] =16'd48;
		memory[665] =16'd26;
		memory[666] =16'd40;
		memory[667] =16'd18;
		memory[668] =16'd21;
		memory[669] =16'd23;
		memory[670] =16'd14;
		memory[671] =16'd42;
		memory[672] =16'd40;
		memory[673] =16'd20;
		memory[674] =16'd11;
		memory[675] =16'd21;
		memory[676] =16'd19;
		memory[677] =16'd30;
		memory[678] =16'd11;
		memory[679] =16'd1;
		memory[680] =16'd37;
		memory[681] =16'd26;
		memory[682] =16'd4;
		memory[683] =16'd29;
		memory[684] =16'd30;
		memory[685] =16'd15;
		memory[686] =16'd6;
		memory[687] =16'd39;
		memory[688] =16'd18;
		memory[689] =16'd3;
		memory[690] =16'd20;
		memory[691] =16'd8;
		memory[692] =16'd0;
		memory[693] =16'd40;
		memory[694] =16'd11;
		memory[695] =16'd36;
		memory[696] =16'd43;
		memory[697] =16'd6;
		memory[698] =16'd1;
		memory[699] =16'd15;
		memory[700] =16'd3;
		memory[701] =16'd38;
		memory[702] =16'd16;
		memory[703] =16'd48;
		memory[704] =16'd27;
		memory[705] =16'd27;
		memory[706] =16'd22;
		memory[707] =16'd45;
		memory[708] =16'd20;
		memory[709] =16'd21;
		memory[710] =16'd31;
		memory[711] =16'd0;
		memory[712] =16'd30;
		memory[713] =16'd24;
		memory[714] =16'd44;
		memory[715] =16'd20;
		memory[716] =16'd34;
		memory[717] =16'd14;
		memory[718] =16'd26;
		memory[719] =16'd38;
		memory[720] =16'd30;
		memory[721] =16'd17;
		memory[722] =16'd13;
		memory[723] =16'd36;
		memory[724] =16'd32;
		memory[725] =16'd11;
		memory[726] =16'd49;
		memory[727] =16'd13;
		memory[728] =16'd49;
		memory[729] =16'd40;
		memory[730] =16'd30;
		memory[731] =16'd0;
		memory[732] =16'd24;
		memory[733] =16'd13;
		memory[734] =16'd7;
		memory[735] =16'd34;
		memory[736] =16'd44;
		memory[737] =16'd40;
		memory[738] =16'd47;
		memory[739] =16'd22;
		memory[740] =16'd47;
		memory[741] =16'd17;
		memory[742] =16'd30;
		memory[743] =16'd19;
		memory[744] =16'd30;
		memory[745] =16'd26;
		memory[746] =16'd40;
		memory[747] =16'd5;
		memory[748] =16'd4;
		memory[749] =16'd13;
		memory[750] =16'd36;
		memory[751] =16'd19;
		memory[752] =16'd7;
		memory[753] =16'd48;
		memory[754] =16'd43;
		memory[755] =16'd20;
		memory[756] =16'd38;
		memory[757] =16'd30;
		memory[758] =16'd44;
		memory[759] =16'd1;
		memory[760] =16'd3;
		memory[761] =16'd43;
		memory[762] =16'd5;
		memory[763] =16'd33;
		memory[764] =16'd16;
		memory[765] =16'd1;
		memory[766] =16'd17;
		memory[767] =16'd48;
		memory[768] =16'd5;
		memory[769] =16'd14;
		memory[770] =16'd5;
		memory[771] =16'd8;
		memory[772] =16'd15;
		memory[773] =16'd48;
		memory[774] =16'd26;
		memory[775] =16'd41;
		memory[776] =16'd20;
		memory[777] =16'd9;
		memory[778] =16'd4;
		memory[779] =16'd34;
		memory[780] =16'd32;
		memory[781] =16'd3;
		memory[782] =16'd36;
		memory[783] =16'd42;
		memory[784] =16'd26;
		memory[785] =16'd27;
		memory[786] =16'd20;
		memory[787] =16'd30;
		memory[788] =16'd16;
		memory[789] =16'd19;
		memory[790] =16'd28;
		memory[791] =16'd22;
		memory[792] =16'd26;
		memory[793] =16'd5;
		memory[794] =16'd1;
		memory[795] =16'd18;
		memory[796] =16'd27;
		memory[797] =16'd37;
		memory[798] =16'd4;
		memory[799] =16'd24;
		memory[800] =16'd47;
		memory[801] =16'd27;
		memory[802] =16'd39;
		memory[803] =16'd10;
		memory[804] =16'd12;
		memory[805] =16'd47;
		memory[806] =16'd26;
		memory[807] =16'd6;
		memory[808] =16'd41;
		memory[809] =16'd47;
		memory[810] =16'd24;
		memory[811] =16'd13;
		memory[812] =16'd21;
		memory[813] =16'd10;
		memory[814] =16'd19;
		memory[815] =16'd16;
		memory[816] =16'd49;
		memory[817] =16'd10;
		memory[818] =16'd46;
		memory[819] =16'd4;
		memory[820] =16'd44;
		memory[821] =16'd46;
		memory[822] =16'd27;
		memory[823] =16'd36;
		memory[824] =16'd41;
		memory[825] =16'd20;
		memory[826] =16'd34;
		memory[827] =16'd27;
		memory[828] =16'd4;
		memory[829] =16'd31;
		memory[830] =16'd29;
		memory[831] =16'd23;
		memory[832] =16'd10;
		memory[833] =16'd31;
		memory[834] =16'd26;
		memory[835] =16'd16;
		memory[836] =16'd14;
		memory[837] =16'd1;
		memory[838] =16'd46;
		memory[839] =16'd18;
		memory[840] =16'd39;
		memory[841] =16'd40;
		memory[842] =16'd7;
		memory[843] =16'd44;
		memory[844] =16'd40;
		memory[845] =16'd37;
		memory[846] =16'd27;
		memory[847] =16'd38;
		memory[848] =16'd7;
		memory[849] =16'd14;
		memory[850] =16'd12;
		memory[851] =16'd42;
		memory[852] =16'd26;
		memory[853] =16'd37;
		memory[854] =16'd3;
		memory[855] =16'd43;
		memory[856] =16'd30;
		memory[857] =16'd6;
		memory[858] =16'd19;
		memory[859] =16'd11;
		memory[860] =16'd17;
		memory[861] =16'd21;
		memory[862] =16'd44;
		memory[863] =16'd35;
		memory[864] =16'd44;
		memory[865] =16'd28;
		memory[866] =16'd43;
		memory[867] =16'd4;
		memory[868] =16'd42;
		memory[869] =16'd47;
		memory[870] =16'd23;
		memory[871] =16'd36;
		memory[872] =16'd45;
		memory[873] =16'd4;
		memory[874] =16'd30;
		memory[875] =16'd37;
		memory[876] =16'd39;
		memory[877] =16'd46;
		memory[878] =16'd39;
		memory[879] =16'd42;
		memory[880] =16'd8;
		memory[881] =16'd28;
		memory[882] =16'd8;
		memory[883] =16'd3;
		memory[884] =16'd40;
		memory[885] =16'd23;
		memory[886] =16'd13;
		memory[887] =16'd8;
		memory[888] =16'd14;
		memory[889] =16'd36;
		memory[890] =16'd41;
		memory[891] =16'd0;
		memory[892] =16'd1;
		memory[893] =16'd15;
		memory[894] =16'd26;
		memory[895] =16'd27;
		memory[896] =16'd9;
		memory[897] =16'd4;
		memory[898] =16'd23;
		memory[899] =16'd18;
		memory[900] =16'd2;
		memory[901] =16'd19;
		memory[902] =16'd15;
		memory[903] =16'd44;

		memory[904] =16'd0;
		memory[905] =16'd0;
		memory[906] =16'd0;
		memory[907] =16'd0;
		memory[908] =16'd0;
		memory[909] =16'd0;
		memory[910] =16'd0;
		memory[911] =16'd0;
		memory[912] =16'd0;
		memory[913] =16'd0;
		memory[914] =16'd0;
		memory[915] =16'd0;
		memory[916] =16'd0;
		memory[917] =16'd0;
		memory[918] =16'd0;
		memory[919] =16'd0;
		memory[920] =16'd0;
		memory[921] =16'd0;
		memory[922] =16'd0;
		memory[923] =16'd0;
		memory[924] =16'd0;
		memory[925] =16'd0;
		memory[926] =16'd0;
		memory[927] =16'd0;
		memory[928] =16'd0;
		memory[929] =16'd0;
		memory[930] =16'd0;
		memory[931] =16'd0;
		memory[932] =16'd0;
		memory[933] =16'd0;
		memory[934] =16'd0;
		memory[935] =16'd0;
		memory[936] =16'd0;
		memory[937] =16'd0;
		memory[938] =16'd0;
		memory[939] =16'd0;
		memory[940] =16'd0;
		memory[941] =16'd0;
		memory[942] =16'd0;
		memory[943] =16'd0;
		memory[944] =16'd0;
		memory[945] =16'd0;
		memory[946] =16'd0;
		memory[947] =16'd0;
		memory[948] =16'd0;
		memory[949] =16'd0;
		memory[950] =16'd0;
		memory[951] =16'd0;
		memory[952] =16'd0;
		memory[953] =16'd0;
		memory[954] =16'd0;
		memory[955] =16'd0;
		memory[956] =16'd0;
		memory[957] =16'd0;
		memory[958] =16'd0;
		memory[959] =16'd0;
		memory[960] =16'd0;
		memory[961] =16'd0;
		memory[962] =16'd0;
		memory[963] =16'd0;
		memory[964] =16'd0;
		memory[965] =16'd0;
		memory[966] =16'd0;
		memory[967] =16'd0;
		memory[968] =16'd0;
		memory[969] =16'd0;
		memory[970] =16'd0;
		memory[971] =16'd0;
		memory[972] =16'd0;
		memory[973] =16'd0;
		memory[974] =16'd0;
		memory[975] =16'd0;
		memory[976] =16'd0;
		memory[977] =16'd0;
		memory[978] =16'd0;
		memory[979] =16'd0;
		memory[980] =16'd0;
		memory[981] =16'd0;
		memory[982] =16'd0;
		memory[983] =16'd0;
		memory[984] =16'd0;
		memory[985] =16'd0;
		memory[986] =16'd0;
		memory[987] =16'd0;
		memory[988] =16'd0;
		memory[989] =16'd0;
		memory[990] =16'd0;
		memory[991] =16'd0;
		memory[992] =16'd0;
		memory[993] =16'd0;
		memory[994] =16'd0;
		memory[995] =16'd0;
		memory[996] =16'd0;
		memory[997] =16'd0;
		memory[998] =16'd0;
		memory[999] =16'd0;
		memory[1000] =16'd0;
		memory[1001] =16'd0;
		memory[1002] =16'd0;
		memory[1003] =16'd0;
		memory[1004] =16'd0;
		memory[1005] =16'd0;
		memory[1006] =16'd0;
		memory[1007] =16'd0;
		memory[1008] =16'd0;
		memory[1009] =16'd0;
		memory[1010] =16'd0;
		memory[1011] =16'd0;
		memory[1012] =16'd0;
		memory[1013] =16'd0;
		memory[1014] =16'd0;
		memory[1015] =16'd0;
		memory[1016] =16'd0;
		memory[1017] =16'd0;
		memory[1018] =16'd0;
		memory[1019] =16'd0;
		memory[1020] =16'd0;
		memory[1021] =16'd0;
		memory[1022] =16'd0;
		memory[1023] =16'd0;
		memory[1024] =16'd0;
		memory[1025] =16'd0;
		memory[1026] =16'd0;
		memory[1027] =16'd0;
		memory[1028] =16'd0;
		memory[1029] =16'd0;
		memory[1030] =16'd0;
		memory[1031] =16'd0;
		memory[1032] =16'd0;
		memory[1033] =16'd0;
		memory[1034] =16'd0;
		memory[1035] =16'd0;
		memory[1036] =16'd0;
		memory[1037] =16'd0;
		memory[1038] =16'd0;
		memory[1039] =16'd0;
		memory[1040] =16'd0;
		memory[1041] =16'd0;
		memory[1042] =16'd0;
		memory[1043] =16'd0;
		memory[1044] =16'd0;
		memory[1045] =16'd0;
		memory[1046] =16'd0;
		memory[1047] =16'd0;
		memory[1048] =16'd0;
		memory[1049] =16'd0;
		memory[1050] =16'd0;
		memory[1051] =16'd0;
		memory[1052] =16'd0;
		memory[1053] =16'd0;
		memory[1054] =16'd0;
		memory[1055] =16'd0;
		memory[1056] =16'd0;
		memory[1057] =16'd0;
		memory[1058] =16'd0;
		memory[1059] =16'd0;
		memory[1060] =16'd0;
		memory[1061] =16'd0;
		memory[1062] =16'd0;
		memory[1063] =16'd0;
		memory[1064] =16'd0;
		memory[1065] =16'd0;
		memory[1066] =16'd0;
		memory[1067] =16'd0;
		memory[1068] =16'd0;
		memory[1069] =16'd0;
		memory[1070] =16'd0;
		memory[1071] =16'd0;
		memory[1072] =16'd0;
		memory[1073] =16'd0;
		memory[1074] =16'd0;
		memory[1075] =16'd0;
		memory[1076] =16'd0;
		memory[1077] =16'd0;
		memory[1078] =16'd0;
		memory[1079] =16'd0;
		memory[1080] =16'd0;
		memory[1081] =16'd0;
		memory[1082] =16'd0;
		memory[1083] =16'd0;
		memory[1084] =16'd0;
		memory[1085] =16'd0;
		memory[1086] =16'd0;
		memory[1087] =16'd0;
		memory[1088] =16'd0;
		memory[1089] =16'd0;
		memory[1090] =16'd0;
		memory[1091] =16'd0;
		memory[1092] =16'd0;
		memory[1093] =16'd0;
		memory[1094] =16'd0;
		memory[1095] =16'd0;
		memory[1096] =16'd0;
		memory[1097] =16'd0;
		memory[1098] =16'd0;
		memory[1099] =16'd0;
		memory[1100] =16'd0;
		memory[1101] =16'd0;
		memory[1102] =16'd0;
		memory[1103] =16'd0;
		memory[1104] =16'd0;
		memory[1105] =16'd0;
		memory[1106] =16'd0;
		memory[1107] =16'd0;
		memory[1108] =16'd0;
		memory[1109] =16'd0;
		memory[1110] =16'd0;
		memory[1111] =16'd0;
		memory[1112] =16'd0;
		memory[1113] =16'd0;
		memory[1114] =16'd0;
		memory[1115] =16'd0;
		memory[1116] =16'd0;
		memory[1117] =16'd0;
		memory[1118] =16'd0;
		memory[1119] =16'd0;
		memory[1120] =16'd0;
		memory[1121] =16'd0;
		memory[1122] =16'd0;
		memory[1123] =16'd0;
		memory[1124] =16'd0;
		memory[1125] =16'd0;
		memory[1126] =16'd0;
		memory[1127] =16'd0;
		memory[1128] =16'd0;
		memory[1129] =16'd0;
		memory[1130] =16'd0;
		memory[1131] =16'd0;
		memory[1132] =16'd0;
		memory[1133] =16'd0;
		memory[1134] =16'd0;
		memory[1135] =16'd0;
		memory[1136] =16'd0;
		memory[1137] =16'd0;
		memory[1138] =16'd0;
		memory[1139] =16'd0;
		memory[1140] =16'd0;
		memory[1141] =16'd0;
		memory[1142] =16'd0;
		memory[1143] =16'd0;
		memory[1144] =16'd0;
		memory[1145] =16'd0;
		memory[1146] =16'd0;
		memory[1147] =16'd0;
		memory[1148] =16'd0;
		memory[1149] =16'd0;
		memory[1150] =16'd0;
		memory[1151] =16'd0;
		memory[1152] =16'd0;
		memory[1153] =16'd0;
		memory[1154] =16'd0;
		memory[1155] =16'd0;
		memory[1156] =16'd0;
		memory[1157] =16'd0;
		memory[1158] =16'd0;
		memory[1159] =16'd0;
		memory[1160] =16'd0;
		memory[1161] =16'd0;
		memory[1162] =16'd0;
		memory[1163] =16'd0;
		memory[1164] =16'd0;
		memory[1165] =16'd0;
		memory[1166] =16'd0;
		memory[1167] =16'd0;
		memory[1168] =16'd0;
		memory[1169] =16'd0;
		memory[1170] =16'd0;
		memory[1171] =16'd0;
		memory[1172] =16'd0;
		memory[1173] =16'd0;
		memory[1174] =16'd0;
		memory[1175] =16'd0;
		memory[1176] =16'd0;
		memory[1177] =16'd0;
		memory[1178] =16'd0;
		memory[1179] =16'd0;
		memory[1180] =16'd0;
		memory[1181] =16'd0;
		memory[1182] =16'd0;
		memory[1183] =16'd0;
		memory[1184] =16'd0;
		memory[1185] =16'd0;
		memory[1186] =16'd0;
		memory[1187] =16'd0;
		memory[1188] =16'd0;
		memory[1189] =16'd0;
		memory[1190] =16'd0;
		memory[1191] =16'd0;
		memory[1192] =16'd0;
		memory[1193] =16'd0;
		memory[1194] =16'd0;
		memory[1195] =16'd0;
		memory[1196] =16'd0;
		memory[1197] =16'd0;
		memory[1198] =16'd0;
		memory[1199] =16'd0;
		memory[1200] =16'd0;
		memory[1201] =16'd0;
		memory[1202] =16'd0;
		memory[1203] =16'd0;
		memory[1204] =16'd0;
		memory[1205] =16'd0;
		memory[1206] =16'd0;
		memory[1207] =16'd0;
end

integer i;
always @(posedge clk) begin
    if(read==1) begin
        for(i=0; i<NO_OF_CORES; i=i+1) begin
             data_out[DATA_LEN*i +: DATA_LEN] <= memory[address[ADDRESS_LEN*i +: ADDRESS_LEN]];
         end
    end
    else if(write==1) begin
         for(i=0; i<NO_OF_CORES; i=i+1) begin
             memory[address[ADDRESS_LEN*i +: ADDRESS_LEN]] <= data_in[DATA_LEN*i +: DATA_LEN];
         end
    end
end
endmodule